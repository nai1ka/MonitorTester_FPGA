module color_lines(


always @(x|y)
begin

end

endmodule